module halfAdder(in1,in2,sum,cout);

input in1,in2;
output sum, cout;
sum=in1^in2;
cout=in1&in2;

endmodule 

 