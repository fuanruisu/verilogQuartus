module Lab3(

	

	//////////// LED //////////
	output		     [9:0]		LEDR,

	//////////// SW //////////
	input 		     [9:0]		SW
);



//=======================================================
//  REG/WIRE declarations
//=======================================================



//=======================================================
//  Structural coding
//=======================================================
 //2-to-1 MUX

assign LEDR[0] = ((~SW[9]&((~SW[8]&SW[0]) | (SW[8]&SW[2]))) | (SW[9]&((~SW[8]&SW[4])|(SW[8]&SW[6]))));
assign LEDR[1] = ((~SW[9]&((~SW[8]&SW[1]) | (SW[8]&SW[3]))) | (SW[9]&((~SW[8]&SW[5])|(SW[8]&SW[7]))));




endmodule
