module Lab2(

	

	//////////// LED //////////
	output		     [3:0]		LEDR,

	//////////// SW //////////
	input 		     [9:0]		SW
);



//=======================================================
//  REG/WIRE declarations
//=======================================================




//=======================================================
//  Structural coding
//=======================================================
 //2-to-1 MUX
assign LEDR[0] = (~SW[9]&SW[0])|(SW[9]&SW[4]);
assign LEDR[1] = (~SW[9]&SW[1])|(SW[9]&SW[5]);
assign LEDR[2] = (~SW[9]&SW[2])|(SW[9]&SW[6]);
assign LEDR[3] = (~SW[9]&SW[3])|(SW[9]&SW[7]);



endmodule
